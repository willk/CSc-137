`include "bcd_mux.v"

module bcd_tester ()
